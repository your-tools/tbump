module test();
    logic [128:0] version_two = "1.2.41-alpha-1";
endmodule
