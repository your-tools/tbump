module test();
    logic [128:0] version = "1.2.41-alpha-1";
endmodule
